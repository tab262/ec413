`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:56:22 11/14/2013 
// Design Name: 
// Module Name:    selectJorBranch 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
/*
module selectJorBranch(
	input[15:0] J_ID_PC,Branch_ID_PC,
	input Branch,selectPCcontrol,
	output[15:0] ID_PC,
	output PCSource);
	
	
	function PCSource, [15:0]f_ID_PC;
		input[15:0] J_ID_PC, Branch_ID_PC;
	if(instruction[31:26] == 6'b000001) begin
		


endmodule
*/